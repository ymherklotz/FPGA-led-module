`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yann Herklotz
// 
// Create Date:    23:10:42 02/19/2017 
// Design Name: 
// Module Name:    led 
// Project Name: 
// Target Devices: Papilio Pro
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module led(
    );


endmodule
